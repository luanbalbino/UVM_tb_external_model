interface mux_if();

  logic [3:0] a,b,c,d;
  logic [1:0] sel;
  logic en;
  logic [3:0] y;

endinterface